// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

#define    d0    D0
#define    d1    D1
#define    d2    D2
#define    d3    D3
#define    d4    D4
#define    d5    D5
#define    d6    D6
#define    d7    D7
#define    d8    D8
#define    rx    RX
#define    tx    TX
#define    a0    A0
#define    sd3   SD3
#define    sd2   SD2
#define    cmd   CMD
#define    sd0   SD0
#define    clk   CLK


fn init() {

}

