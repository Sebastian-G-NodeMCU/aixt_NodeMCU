// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pwm.c.v
// Author: Fernando Martínez Santa - Sebastian Gongora  - Brayan Gaitan
// Date: 2024
// License: MIT
//
// // Description: PWM functions (Ai_Thinker_Ai-WB2-32S-Kit)

module pwm

fn init() {

}